//-----------------------------------------------------
// PROYECTO 1  : SD HOST
// Archivo     : testfisico.v
// Descripcion : testbench para capa física de bloque de DATA
// Estudiante  : Mario Castresana Avendaño - A41267
//-----------------------------------------------------

`timescale 1ns / 1ps

//`include "DATA.v"
`include "probador.v"
`include "DATA_PHYSICAL.v"




module testbench;


// Wires para probar data


//salidas de capa física
 
      
//probador para bloque de control de datos
probador DataTest(


);

// Instanciar Unit Under Test (UUT) DATA
DATA DATA_CONTROL(
	//inputs

	//outputs
      
);

endmodule