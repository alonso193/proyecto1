//el siguiente módulo se encarga de la transferencia de comandos del sdHost a la sdCard y de la sdCard hacia el sdHost
module CMD (input clk, reset);

endmodule // CMD
